`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/05/2023 03:36:42 PM
// Design Name: 
// Module Name: TapeStorage
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TapeStorage( input clk, BlockRamConnection.owner stringRam, BlockRamConnection.owner structRam);
    BlockRamSharer #(.NUMWORDS(Core::StringTapeLength)) stringTapeRam (.clk, .r(stringRam));
    BlockRamSharer #(.NUMWORDS(Core::StructTapeLength)) structTapeRam (.clk, .r(structRam));
endmodule
